                                                                                ░░░░░░░░░░░█▀▀░░█░░░░░░
                                                                                ░░░░░░▄▀▀▀▀░░░░░█▄▄░░░░
                                                                                ░░░░░░█░█░░░░░░░░░░▐░░░
                                                                                ░░░░░░▐▐░░░░░░░░░▄░▐░░░
                                                                                ░░░░░░█░░░░░░░░▄▀▀░▐░░░
                                                                                ░░░░▄▀░░░░░░░░▐░▄▄▀░░░░
                                                                                ░░▄▀░░░▐░░░░░█▄▀░▐░░░░░
                                                                                ░░█░░░▐░░░░░░░░▄░█░░░░░
                                                                                ░░░█▄░░▀▄░░░░▄▀▐░█░░░░░
                                                                                ░░░█▐▀▀▀░▀▀▀▀░░▐░█░░░░░
                                                                                ░░▐█▐▄░░▀░░░░░░▐░█▄▄░░
                                                                                ░░░▀▀░▄TSM▄░░░▐▄▄▄▀░░░

                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢰⣶⡄⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢀⣀⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢴⣄⡀⠀⠀⠀⠀⠀⠀⠀⢈⣧⣷⡤⠄⠀⠀⠀⠀⠀⠀⢠⣄⡀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⠀⢀⣾⡿⠛⠃⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠸⣿⣄⠀⠀⠀⠀⠀⠀⠀⠀⣽⣿⠀⠀⠀⠀⠀⠀⠀⠀⠀⠻⣷⡀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠰⠤⣶⡷⢢⡀⠀⠀⠀⢸⣿⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢈⣿⡅⠀⠀⠀⢀⣴⡿⠟⠛⠋⠀⠀⠀⠀⢀⣄⠀⠀⠀⠀⢹⡇⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠉⠉⠁⠀⠀⠀⠈⣿⣧⠄⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢰⡿⠋⠀⠀⠀⠀⢹⣿⠁⠀⠀⠀⠀⠀⠀⠀⢸⣿⠀⠀⠀⢀⣼⡇⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠘⣿⡆⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢸⡄⠀⠀⠀⠀⠀⠘⣿⣆⠀⠀⠀⠀⠀⠀⣴⣿⠏⠀⠀⣰⡿⠋⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⡀⠀⠀⠘⣿⣆⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠉⢿⡄⠂⠀⠀⠀⠀⢈⣿⡇⠀⠀⠀⠀⠸⣿⡀⠀⠀⠸⣿⠤⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⣀⠞⠀⠀⠀⠀⠸⣿⠀⠀⠀⠀⠀⠀⠀⠑⣄⡀⠀⠀⠀⠀⢻⠀⠀⠀⠀⢴⡟⠋⠀⠀⠀⠀⠀⠀⠹⣿⣜⠁⠀⠙⠷⣄⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠈⣿⠀⠀⠀⠀⠀⣸⡟⠀⠀⠀⠀⠀⠀⠀⠀⢠⣉⡀⠀⠐⠒⠚⠁⠠⠄⠀⢸⣦⠄⠀⠀⠐⠀⠀⠀⠀⠈⢿⡆⠀⠀⠀⢸⡇⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⢠⡿⠀⠀⠀⢀⣼⠋⠀⠀⠀⠀⠀⠀⠀⠀⠀⣸⠉⣿⠀⠀⠀⠀⠀⠀⠀⠀⠈⢿⡄⠀⠀⠀⠀⠀⠀⢀⣴⡟⠁⠀⠀⠀⠀⠀⢀⣀⣀⣦⠀⠀⡄
                                                    ⠀⠀⠀⠀⢀⡟⠁⠀⠀⠀⢸⠃⠀⠀⠀⠀⠀⠀⠀⠀⢀⣼⠏⠀⢿⡄⠀⠀⠀⠀⠀⠀⠀⠀⣸⠇⠀⠀⠀⠀⠀⣴⡟⠁⠀⠀⠀⠀⠀⠀⠀⠘⠶⠖⠛⠈⠉⠀
                                                    ⠀⠀⠀⠀⢸⠀⠀⠀⠀⠀⣹⠀⠀⠀⠀⠀⠀⢀⣤⡾⠟⠁⠀⠀⠈⠻⢶⣤⣀⣀⠀⠀⠀⠊⠁⠀⠀⠀⠀⠀⠀⣿⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠸⡀⠀⠀⠀⠀⠸⡇⠀⠀⠀⠀⢀⣿⠋⠀⠀⠀⠀⢄⣰⠲⡤⡀⠌⠛⢷⣄⠀⠀⠀⠀⠀⠀⠀⠀⠀⠈⠻⣦⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠁⠀⠀⠀⠀⠀⠉⠀⠀⠀⠀⢸⡏⠐⡂⠐⠀⠀⠀⠈⠙⠒⠲⠤⠤⠾⠟⠛⢻⢷⣦⣀⠀⠀⠀⠀⠀⠀⠈⣧⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠘⣷⡀⠃⠀⠀⡄⠀⠀⠀⠀⢤⠂⠀⠐⠀⢧⡈⠀⢯⡻⣷⡀⠀⠀⠀⠀⠀⠋⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢀⣠⣽⣷⣄⠀⠀⠃⠳⠸⡄⠄⠀⠀⠀⠀⠀⢀⣀⢀⠀⣅⢸⣿⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢀⣠⡾⠟⠉⠀⣨⠙⠛⠶⠤⣀⣀⠀⠀⠀⠀⠰⠤⢣⢸⡘⣌⡆⠘⠀⣿⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢠⡿⣫⡀⠀⢠⠖⡇⠀⠀⡀⠀⠀⠀⠀⠀⢀⣀⠀⠀⠠⠤⣅⣈⣠⣴⢾⣿⣀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢠⣿⠑⣿⣡⠤⡏⣠⢯⠀⠊⠁⡀⠀⠀⠀⠀⠈⠉⡟⠛⠐⠰⠀⠀⠇⢷⡀⠟⠛⠻⣶⣤⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠘⣿⣼⡵⠃⢰⠃⢀⡞⢠⠀⠀⠇⠀⠀⠀⠀⣰⠶⠃⠀⠀⠀⠀⠀⠀⠀⠹⣄⠀⢄⠲⠙⢿⣆⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⠀⠀⣠⣶⡿⠟⠉⠀⠀⠁⠀⠈⠀⠈⠀⢠⡶⣆⠀⠀⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠘⡆⠸⣤⡘⠈⣿⡄⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠀⣠⣾⠟⣥⢰⠆⢠⣄⠀⠀⠀⢀⡀⠀⠀⠘⠁⠙⠀⠀⠁⠀⠀⠀⠀⠀⢀⠀⢤⠘⡆⠸⣄⢳⠀⣇⣹⣶⣿⣧⣀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⣰⣿⠃⠰⠃⠚⠀⠈⠁⠽⠄⠀⠀⠉⠙⠒⠦⠤⣄⣀⣀⣀⣀⣀⣀⣀⢀⣘⣂⣘⣃⣷⣤⣽⡾⠿⠟⠛⣉⢈⠙⣿⣧⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⢀⣿⠇⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⣀⠀⠀⠀⠀⠀⠀⠈⣍⣉⢉⠉⠛⠛⠛⠛⠋⠉⠉⠉⠀⠀⠀⠀⠀⠹⡌⠂⠁⢻⣷⡀⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⢸⣿⠀⢷⣆⡀⠀⠀⠀⠀⠀⠀⠀⠀⠉⢠⠀⠀⠀⠀⠀⠀⠈⠛⠎⠃⠀⠀⠀⠀⢠⠀⣄⠀⡦⠀⢰⠀⠀⡀⢀⠰⡶⡄⣿⡇⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠸⣿⡀⠘⢸⢹⣆⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⡀⠄⠀⠀⠀⠀⢠⡀⣤⢰⡆⣸⠀⣿⠀⠷⠀⠈⡀⣌⢿⠈⡇⠇⠁⣿⡇⠀⠀⠀⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⠀⠻⣷⡄⠘⠼⢸⠁⡇⢰⠀⡄⠀⠀⠀⡴⠀⠀⠰⠃⠀⠀⠀⠀⠀⠀⠟⠓⠺⠃⢙⠀⢁⡀⣤⢇⠀⢣⢸⡸⡆⠟⢀⣼⡿⠁⡴⠀⣄⠀⠀⠀⠀⠀
                                                    ⠀⠀⠀⠀⢀⣠⣿⣿⣄⠀⡄⣤⡀⠈⡄⢀⡀⠀⠀⠃⠸⠰⠃⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠈⡇⠘⠂⠛⠸⠄⠘⠋⠁⣠⣤⣾⠟⢡⠞⢁⡴⠋⢰⡄⠀⠀⠀
                                                    ⠀⠀⠀⠶⣫⠵⠋⣩⢿⣷⣝⣁⡇⢀⠇⢸⠀⡆⢠⡀⢰⠀⡀⠀⠀⠀⢠⡀⡄⣦⠠⡄⠒⠒⠀⠀⠀⠀⠀⢀⣠⣤⣶⡿⢟⡿⢁⡴⠋⣠⠞⠁⣠⠞⠁⠀⠀⠀
                                                    ⠀⠀⠐⣋⣡⠖⠋⠁⣠⠼⠛⠿⢿⣶⣶⣬⣄⣃⣈⣀⣈⣀⠀⠀⠀⠀⠀⢀⣈⣙⣀⣀⣀⣤⣤⣶⣶⣾⠿⠿⢛⡿⠁⡴⠋⣠⠎⢀⡾⠃⢀⣴⠃⠀⠴⠀⠀⠀
