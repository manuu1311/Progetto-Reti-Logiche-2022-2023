                                                                                ░░░░░░░░░░░█▀▀░░█░░░░░░
                                                                                ░░░░░░▄▀▀▀▀░░░░░█▄▄░░░░
                                                                                ░░░░░░█░█░░░░░░░░░░▐░░░
                                                                                ░░░░░░▐▐░░░░░░░░░▄░▐░░░
                                                                                ░░░░░░█░░░░░░░░▄▀▀░▐░░░
                                                                                ░░░░▄▀░░░░░░░░▐░▄▄▀░░░░
                                                                                ░░▄▀░░░▐░░░░░█▄▀░▐░░░░░
                                                                                ░░█░░░▐░░░░░░░░▄░█░░░░░
                                                                                ░░░█▄░░▀▄░░░░▄▀▐░█░░░░░
                                                                                ░░░█▐▀▀▀░▀▀▀▀░░▐░█░░░░░
                                                                                ░░▐█▐▄░░▀░░░░░░▐░█▄▄░░
                                                                                ░░░▀▀░▄    ▄░░░▐▄▄▄▀░░░                                         
                                                                                  
                                                                                  
                                                                                  
                                                                                  
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢰⣶⡄⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢀⣀⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢴⣄⡀⠀⠀⠀⠀⠀⠀⠀⢈⣧⣷⡤⠄⠀⠀⠀⠀⠀⠀⢠⣄⡀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⢀⣾⡿⠛⠃⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠸⣿⣄⠀⠀⠀⠀⠀⠀⠀⠀⣽⣿⠀⠀⠀⠀⠀⠀⠀⠀⠀⠻⣷⡀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠰⠤⣶⡷⢢⡀⠀⠀⠀⢸⣿⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢈⣿⡅⠀⠀⠀⢀⣴⡿⠟⠛⠋⠀⠀⠀⠀⢀⣄⠀⠀⠀⠀⢹⡇⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠉⠉⠁⠀⠀⠀⠈⣿⣧⠄⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢰⡿⠋⠀⠀⠀⠀⢹⣿⠁⠀⠀⠀⠀⠀⠀⠀⢸⣿⠀⠀⠀⢀⣼⡇⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠘⣿⡆⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢸⡄⠀⠀⠀⠀⠀⠘⣿⣆⠀⠀⠀⠀⠀⠀⣴⣿⠏⠀⠀⣰⡿⠋⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⡀⠀⠀⠘⣿⣆⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠉⢿⡄⠂⠀⠀⠀⠀⢈⣿⡇⠀⠀⠀⠀⠸⣿⡀⠀⠀⠸⣿⠤⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⣀⠞⠀⠀⠀⠀⠸⣿⠀⠀⠀⠀⠀⠀⠀⠑⣄⡀⠀⠀⠀⠀⢻⠀⠀⠀⠀⢴⡟⠋⠀⠀⠀⠀⠀⠀⠹⣿⣜⠁⠀⠙⠷⣄⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠈⣿⠀⠀⠀⠀⠀⣸⡟⠀⠀⠀⠀⠀⠀⠀⠀⢠⣉⡀⠀⠐⠒⠚⠁⠠⠄⠀⢸⣦⠄⠀⠀⠐⠀⠀⠀⠀⠈⢿⡆⠀⠀⠀⢸⡇⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⢠⡿⠀⠀⠀⢀⣼⠋⠀⠀⠀⠀⠀⠀⠀⠀⠀⣸⠉⣿⠀⠀⠀⠀⠀⠀⠀⠀⠈⢿⡄⠀⠀⠀⠀⠀⠀⢀⣴⡟⠁⠀⠀⠀⠀⠀⢀⣀⣀⣦⠀⠀⡄
                                                      ⠀⠀⠀⠀⢀⡟⠁⠀⠀⠀⢸⠃⠀⠀⠀⠀⠀⠀⠀⠀⢀⣼⠏⠀⢿⡄⠀⠀⠀⠀⠀⠀⠀⠀⣸⠇⠀⠀⠀⠀⠀⣴⡟⠁⠀⠀⠀⠀⠀⠀⠀⠘⠶⠖⠛⠈⠉⠀
                                                      ⠀⠀⠀⠀⢸⠀⠀⠀⠀⠀⣹⠀⠀⠀⠀⠀⠀⢀⣤⡾⠟⠁⠀⠀⠈⠻⢶⣤⣀⣀⠀⠀⠀⠊⠁⠀⠀⠀⠀⠀⠀⣿⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠸⡀⠀⠀⠀⠀⠸⡇⠀⠀⠀⠀⢀⣿⠋⠀⠀⠀⠀⢄⣰⠲⡤⡀⠌⠛⢷⣄⠀⠀⠀⠀⠀⠀⠀⠀⠀⠈⠻⣦⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠁⠀⠀⠀⠀⠀⠉⠀⠀⠀⠀⢸⡏⠐⡂⠐⠀⠀⠀⠈⠙⠒⠲⠤⠤⠾⠟⠛⢻⢷⣦⣀⠀⠀⠀⠀⠀⠀⠈⣧⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠘⣷⡀⠃⠀⠀⡄⠀⠀⠀⠀⢤⠂⠀⠐⠀⢧⡈⠀⢯⡻⣷⡀⠀⠀⠀⠀⠀⠋⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢀⣠⣽⣷⣄⠀⠀⠃⠳⠸⡄⠄⠀⠀⠀⠀⠀⢀⣀⢀⠀⣅⢸⣿⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢀⣠⡾⠟⠉⠀⣨⠙⠛⠶⠤⣀⣀⠀⠀⠀⠀⠰⠤⢣⢸⡘⣌⡆⠘⠀⣿⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢠⡿⣫⡀⠀⢠⠖⡇⠀⠀⡀⠀⠀⠀⠀⠀⢀⣀⠀⠀⠠⠤⣅⣈⣠⣴⢾⣿⣀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⢠⣿⠑⣿⣡⠤⡏⣠⢯⠀⠊⠁⡀⠀⠀⠀⠀⠈⠉⡟⠛⠐⠰⠀⠀⠇⢷⡀⠟⠛⠻⣶⣤⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠘⣿⣼⡵⠃⢰⠃⢀⡞⢠⠀⠀⠇⠀⠀⠀⠀⣰⠶⠃⠀⠀⠀⠀⠀⠀⠀⠹⣄⠀⢄⠲⠙⢿⣆⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⣠⣶⡿⠟⠉⠀⠀⠁⠀⠈⠀⠈⠀⢠⡶⣆⠀⠀⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠘⡆⠸⣤⡘⠈⣿⡄⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⣠⣾⠟⣥⢰⠆⢠⣄⠀⠀⠀⢀⡀⠀⠀⠘⠁⠙⠀⠀⠁⠀⠀⠀⠀⠀⢀⠀⢤⠘⡆⠸⣄⢳⠀⣇⣹⣶⣿⣧⣀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⣰⣿⠃⠰⠃⠚⠀⠈⠁⠽⠄⠀⠀⠉⠙⠒⠦⠤⣄⣀⣀⣀⣀⣀⣀⣀⢀⣘⣂⣘⣃⣷⣤⣽⡾⠿⠟⠛⣉⢈⠙⣿⣧⡀⠀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⢀⣿⠇⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⣀⠀⠀⠀⠀⠀⠀⠈⣍⣉⢉⠉⠛⠛⠛⠛⠋⠉⠉⠉⠀⠀⠀⠀⠀⠹⡌⠂⠁⢻⣷⡀⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⢸⣿⠀⢷⣆⡀⠀⠀⠀⠀⠀⠀⠀⠀⠉⢠⠀⠀⠀⠀⠀⠀⠈⠛⠎⠃⠀⠀⠀⠀⢠⠀⣄⠀⡦⠀⢰⠀⠀⡀⢀⠰⡶⡄⣿⡇⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠸⣿⡀⠘⢸⢹⣆⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⡀⠄⠀⠀⠀⠀⢠⡀⣤⢰⡆⣸⠀⣿⠀⠷⠀⠈⡀⣌⢿⠈⡇⠇⠁⣿⡇⠀⠀⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠻⣷⡄⠘⠼⢸⠁⡇⢰⠀⡄⠀⠀⠀⡴⠀⠀⠰⠃⠀⠀⠀⠀⠀⠀⠟⠓⠺⠃⢙⠀⢁⡀⣤⢇⠀⢣⢸⡸⡆⠟⢀⣼⡿⠁⡴⠀⣄⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⢀⣠⣿⣿⣄⠀⡄⣤⡀⠈⡄⢀⡀⠀⠀⠃⠸⠰⠃⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠈⡇⠘⠂⠛⠸⠄⠘⠋⠁⣠⣤⣾⠟⢡⠞⢁⡴⠋⢰⡄⠀⠀⠀
                                                      ⠀⠀⠀⠶⣫⠵⠋⣩⢿⣷⣝⣁⡇⢀⠇⢸⠀⡆⢠⡀⢰⠀⡀⠀⠀⠀⢠⡀⡄⣦⠠⡄⠒⠒⠀⠀⠀⠀⠀⢀⣠⣤⣶⡿⢟⡿⢁⡴⠋⣠⠞⠁⣠⠞⠁⠀⠀⠀
                                                      ⠀⠀⠐⣋⣡⠖⠋⠁⣠⠼⠛⠿⢿⣶⣶⣬⣄⣃⣈⣀⣈⣀⠀⠀⠀⠀⠀⢀⣈⣙⣀⣀⣀⣤⣤⣶⣶⣾⠿⠿⢛⡿⠁⡴⠋⣠⠎⢀⡾⠃⢀⣴⠃⠀⠴⠀⠀⠀
                                                      ⠀⠀⠰⠋⠀⢠⠴⠋⠁⠀⣀⡴⠋⠁⣨⠟⠉⣻⠿⠛⣻⠟⠛⣿⠿⠟⢻⠟⠛⢛⡿⠛⣻⠟⠉⠀⣰⠃⢀⡼⠋⠀⠘⠁⠼⠃⠠⠏⠀⠀⠘⠁⠀⠀⠀⠀⠀⠀
                                                      ⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠉⣀⠀⠚⠁⠀⠐⠃⠀⠐⠁⠀⠀⠁⠀⠀⠀⠀⠀⠁⠀⠀⠁⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀⠀
